`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:10:28 04/10/2017 
// Design Name: 
// Module Name:    MUX4T1_5 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module   MUX4T1_5(input [1:0]s,
						 input [4:0]I0,
						 input [4:0]I1,
						 input [4:0]I2,
						 input [4:0]I3,						
						 output reg[4:0]o
						 );

		always @ *//5λ4ѡһ,I0��I1��I2��I3��Ӧѡ��ͨ��0��1��2��3
			case(s)
				2'd0: o <= I0;
				2'd1: o <= I1;
				2'd2: o <= I2;
				2'd3: o <= I3;
			endcase	
endmodule
